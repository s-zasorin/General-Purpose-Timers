module encoder_mode (
  input  logic clk_i    ,
  input  logic aresetn_i,
  input  logic ti1f_i   ,
  input  logic ti2f_i   ,

  output logic clk_1d2_o,
  output logic clk_2d1_o 
);

endmodule